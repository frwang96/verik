`timescale 1ns / 1ns

module Minimal;

endmodule: Minimal