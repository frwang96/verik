module minimal;
    timeunit 1ns / 1ns;

endmodule: minimal