/*
 * SPDX-License-Identifier: Apache-2.0
 */

// test.sv /////////////////////////////////////////////////////////////////////////////////////////////////////////////

typedef enum { E0, E1, E2 } e0;

e0 x0;

class c;

    typedef enum { E3, E4 } e1;

    e1 x1;

endclass
