typedef enum logic [1:0] {
    State_OPENED  = 2'h0,
    State_OPENING = 2'h1,
    State_CLOSED  = 2'h2,
    State_CLOSING = 2'h3
} State;
