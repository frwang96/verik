/*
 * SPDX-License-Identifier: Apache-2.0
 */

// test.sv /////////////////////////////////////////////////////////////////////////////////////////////////////////////

typedef logic [7:0] t0;

t0 x0;

typedef logic t1 [$];

t1 x1;

class c;

    typedef logic t2;

    t2 x2;

endclass
