`timescale 1ns / 1ns

module minimal;

endmodule: minimal