`timescale 1ns / 1ns

package pkg;

    `include "lock.svh"

endpackage
