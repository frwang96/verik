package pkg;
    timeunit 1ns / 1ns;

    `include "lock.svh"
endpackage
