`timescale 1ns / 1ns

package pkg;

    `include "Lock.svh"

endpackage
