/*
 * SPDX-License-Identifier: Apache-2.0
 */

// test.sv /////////////////////////////////////////////////////////////////////////////////////////////////////////////

class c0;
endclass

class c1 extends c0;
endclass

class c2 #(type T, type U, int V = 0);
endclass
