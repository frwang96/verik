typedef enum logic [1:0] {
    STATE_OPENED  = 2'h0,
    STATE_OPENING = 2'h1,
    STATE_CLOSED  = 2'h2,
    STATE_CLOSING = 2'h3
} state;
