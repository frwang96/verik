typedef enum {
    State_OPENED,
    State_OPENING,
    State_CLOSED,
    State_CLOSING
} State;
