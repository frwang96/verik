/*
 * Copyright (c) 2022 Francis Wang
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

// test.sv /////////////////////////////////////////////////////////////////////////////////////////////////////////////

module m0;
endmodule

module m1(
    input logic x0,
    input logic [7:0] x1,
    output logic [3:0][1:0] x2
);
endmodule

module m2(x3, x4);
    input x3;
    input [7:0] x4;
endmodule
