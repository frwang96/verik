package dut_pkg;
    timeunit 1ns / 1ns;

    `include "multiplier.svh"
endpackage
