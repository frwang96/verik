int WIDTH = 8;
