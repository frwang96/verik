`timescale 1ns / 1ns

package dut_pkg;

    `include "multiplier.svh"

endpackage
