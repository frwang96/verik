/*
 * SPDX-License-Identifier: Apache-2.0
 */

// Test0.sv ////////////////////////////////////////////////////////////////////////////////////////////////////////////

module M0;

    M1 m0 (
        .C  ( 8'h00 ),
        .x0 ( 1'b0 ),
        .x1 ( 4'b0000 ),
        .x2 (  )
    );

    M1 m1 (
        .C  ( 8'h00 ),
        .x0 ( 1'b0 ),
        .x1 ( 4'b0000 ),
        .x2 (  )
    );

endmodule : M0

// Test1.sv ////////////////////////////////////////////////////////////////////////////////////////////////////////////

module M1(
    input  logic [7:0] C,
    input  logic       x0,
    input  logic [3:0] x1,
    output logic       x2
);

endmodule : M1
