/*
 * SPDX-License-Identifier: Apache-2.0
 */

// test.sv /////////////////////////////////////////////////////////////////////////////////////////////////////////////

typedef logic [3:0] t;

typedef struct {
    int x0;
    time x1;
    t x2;
} s;

s x3;
