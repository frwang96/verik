/*
 * SPDX-License-Identifier: Apache-2.0
 */

// test.sv /////////////////////////////////////////////////////////////////////////////////////////////////////////////

int x0 [$];

int x1 [string];

logic [3:0][7:0] x3 [1:0];
