/*
 * Copyright (c) 2022 Francis Wang
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

// M.sv ////////////////////////////////////////////////////////////////////////////////////////////////////////////////

`ifndef VERIK
`define VERIK
`timescale 1ns / 1ns
`endif

module M;

    N n1 (
        .A ( 8'h00 ),
        .x ( 1'b0 ),
        .y ( 4'b0000 ),
        .z ( )
    );

    N n2 (
        .A ( 8'h00 ),
        .x ( 1'b0 ),
        .y ( 4'b0000 ),
        .z ( )
    );

endmodule : M

module N(
    input  logic [7:0] A,
    input  logic       x,
    input  logic [3:0] y,
    output logic       z
);

endmodule : N
